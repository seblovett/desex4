magic
tech c035u
timestamp 1387283479
<< pwell >>
rect 9360 0 9560 48
<< metal1 >>
rect 4141 918 4943 928
rect 1861 895 2015 907
rect 4645 896 4799 906
rect 6925 902 9570 912
rect 0 874 4272 884
rect 4286 874 4750 884
rect 4837 874 4991 884
rect 6085 875 6239 885
rect 8293 880 8447 890
rect 0 853 1487 863
rect 1501 852 1967 862
rect 2053 852 2159 862
rect 2245 852 2375 862
rect 2941 854 3071 864
rect 3109 854 3240 864
rect 3661 852 3791 862
rect 3853 852 3935 862
rect 4021 852 5567 862
rect 5581 852 5711 862
rect 5725 852 6191 862
rect 7069 860 7199 870
rect 7789 857 7919 867
rect 7933 857 8399 867
rect 9133 855 9570 865
<< m2contact >>
rect 4127 916 4141 930
rect 4943 916 4957 930
rect 1847 894 1861 908
rect 2015 894 2029 908
rect 4631 894 4645 908
rect 4799 894 4813 908
rect 6911 901 6925 915
rect 4272 872 4286 886
rect 4750 872 4764 886
rect 4823 872 4837 886
rect 4991 872 5005 886
rect 6071 873 6085 887
rect 6239 873 6253 887
rect 8279 878 8293 892
rect 8447 878 8461 892
rect 1487 850 1501 864
rect 1967 850 1981 864
rect 2039 850 2053 864
rect 2159 850 2173 864
rect 2231 850 2245 864
rect 2375 850 2389 864
rect 2927 850 2941 864
rect 3071 850 3085 864
rect 3095 850 3109 864
rect 3240 850 3254 864
rect 3647 850 3661 864
rect 3791 850 3805 864
rect 3839 850 3853 864
rect 3935 850 3949 864
rect 4007 850 4021 864
rect 5567 850 5581 864
rect 5711 850 5725 864
rect 6191 850 6205 864
rect 7055 857 7069 871
rect 7199 858 7213 872
rect 7775 855 7789 869
rect 7919 855 7933 869
rect 8399 855 8413 869
rect 9119 851 9133 865
<< metal2 >>
rect 1536 851 1644 863
rect 1488 847 1500 850
rect 1536 847 1548 851
rect 1632 847 1644 851
rect 1800 847 1812 960
rect 1848 847 1860 894
rect 1944 847 1956 960
rect 1968 847 1980 850
rect 2016 847 2028 894
rect 2040 847 2052 850
rect 2136 847 2148 960
rect 2160 847 2172 850
rect 2208 847 2220 960
rect 2232 847 2244 850
rect 2376 847 2388 850
rect 2928 847 2940 850
rect 3000 847 3012 960
rect 3024 847 3036 960
rect 3072 847 3084 850
rect 3096 847 3108 850
rect 3240 847 3252 850
rect 3648 847 3660 850
rect 3792 847 3804 850
rect 3840 847 3852 850
rect 3936 847 3948 850
rect 4008 847 4020 850
rect 4128 847 4140 916
rect 4200 847 4212 960
rect 4272 847 4284 872
rect 4320 853 4428 865
rect 4320 847 4332 853
rect 4416 847 4428 853
rect 4584 847 4596 960
rect 4632 847 4644 894
rect 4728 847 4740 960
rect 4752 847 4764 872
rect 4800 847 4812 894
rect 4824 847 4836 872
rect 4920 847 4932 960
rect 4944 847 4956 916
rect 4992 847 5004 872
rect 5016 851 5172 863
rect 5016 847 5028 851
rect 5160 847 5172 851
rect 5568 847 5581 850
rect 5712 847 5725 850
rect 5760 851 5868 863
rect 5760 847 5772 851
rect 5856 847 5868 851
rect 6024 847 6036 960
rect 6072 847 6084 873
rect 6168 847 6180 960
rect 6192 847 6204 850
rect 6240 847 6252 873
rect 6264 851 6348 863
rect 6264 847 6276 851
rect 6336 847 6348 851
rect 6384 847 6396 960
rect 6912 847 6924 901
rect 7056 847 7068 857
rect 7128 847 7140 960
rect 7152 847 7164 960
rect 7200 847 7212 858
rect 7224 853 7380 865
rect 7224 847 7236 853
rect 7368 847 7380 853
rect 7776 847 7788 855
rect 7920 847 7932 855
rect 7968 854 8076 866
rect 7968 847 7980 854
rect 8064 847 8076 854
rect 8232 847 8244 960
rect 8280 847 8292 878
rect 8376 847 8388 960
rect 8400 847 8412 855
rect 8448 847 8460 878
rect 8472 856 8556 868
rect 8472 847 8484 856
rect 8544 847 8556 856
rect 8592 847 8604 960
rect 9120 847 9132 851
rect 9360 847 9560 960
rect 0 0 200 48
rect 216 0 228 48
rect 240 0 252 48
rect 264 0 276 48
rect 288 0 300 48
rect 1656 0 1668 48
rect 2784 0 2796 48
rect 3648 0 3660 48
rect 4056 0 4068 48
rect 4440 0 4452 48
rect 5880 0 5892 48
rect 8088 0 8100 48
rect 9360 0 9560 48
use leftbuf leftbuf_0
timestamp 1386242881
transform 1 0 0 0 1 48
box 0 0 1464 799
use inv inv_0
timestamp 1386238110
transform 1 0 1464 0 1 48
box 0 0 120 799
use halfadder halfadder_0
timestamp 1386235204
transform 1 0 1584 0 1 48
box 0 0 312 799
use mux2 mux2_0
timestamp 1386235218
transform 1 0 1896 0 1 48
box 0 0 192 799
use mux2 mux2_1
timestamp 1386235218
transform 1 0 2088 0 1 48
box 0 0 192 799
use scandtype scandtype_0
timestamp 1386241841
transform 1 0 2280 0 1 48
box 0 0 624 799
use tielow tielow_0
timestamp 1386086605
transform 1 0 2904 0 1 48
box 0 0 48 799
use mux2 mux2_2
timestamp 1386235218
transform 1 0 2952 0 1 48
box 0 0 192 799
use scandtype scandtype_1
timestamp 1386241841
transform 1 0 3144 0 1 48
box 0 0 624 799
use inv inv_4
timestamp 1386238110
transform 1 0 3768 0 1 48
box 0 0 120 799
use fulladder fulladder_0
timestamp 1386234928
transform 1 0 3888 0 1 48
box 0 0 360 799
use inv inv_1
timestamp 1386238110
transform 1 0 4248 0 1 48
box 0 0 120 799
use halfadder halfadder_1
timestamp 1386235204
transform 1 0 4368 0 1 48
box 0 0 312 799
use mux2 mux2_3
timestamp 1386235218
transform 1 0 4680 0 1 48
box 0 0 192 799
use mux2 mux2_4
timestamp 1386235218
transform 1 0 4872 0 1 48
box 0 0 192 799
use scandtype scandtype_2
timestamp 1386241841
transform 1 0 5064 0 1 48
box 0 0 624 799
use inv inv_2
timestamp 1386238110
transform 1 0 5688 0 1 48
box 0 0 120 799
use halfadder halfadder_2
timestamp 1386235204
transform 1 0 5808 0 1 48
box 0 0 312 799
use mux2 mux2_5
timestamp 1386235218
transform 1 0 6120 0 1 48
box 0 0 192 799
use scanreg scanreg_0
timestamp 1386241447
transform 1 0 6312 0 1 48
box 0 0 720 799
use tielow tielow_1
timestamp 1386086605
transform 1 0 7032 0 1 48
box 0 0 48 799
use mux2 mux2_6
timestamp 1386235218
transform 1 0 7080 0 1 48
box 0 0 192 799
use scandtype scandtype_4
timestamp 1386241841
transform 1 0 7272 0 1 48
box 0 0 624 799
use inv inv_3
timestamp 1386238110
transform 1 0 7896 0 1 48
box 0 0 120 799
use halfadder halfadder_3
timestamp 1386235204
transform 1 0 8016 0 1 48
box 0 0 312 799
use mux2 mux2_7
timestamp 1386235218
transform 1 0 8328 0 1 48
box 0 0 192 799
use scanreg scanreg_1
timestamp 1386241447
transform 1 0 8520 0 1 48
box 0 0 720 799
use rightend rightend_0
timestamp 1386235834
transform 1 0 9240 0 1 48
box 0 0 320 799
<< labels >>
rlabel metal1 0 853 0 863 3 Operand2
rlabel metal1 0 874 0 884 4 Operand1
rlabel metal2 1656 0 1668 0 1 OP2_INV_Cin
rlabel metal2 4440 0 4452 0 1 OP1_INV_Cin
rlabel metal2 2784 0 2796 0 1 DIVH_1
rlabel metal2 3648 0 3660 0 1 DIVL_1
rlabel metal2 4056 0 4068 0 1 ACC_Cin
rlabel metal2 8088 0 8100 0 1 RESULT_INV_Cin
rlabel metal2 1800 960 1812 960 5 OP2_INV_Cout
rlabel metal2 3024 960 3036 960 5 DIVL_P
rlabel metal2 3000 960 3012 960 5 LOAD_DIVL
rlabel metal2 4584 960 4596 960 1 OP1_INV_Cout
rlabel metal2 4728 960 4740 960 5 INV_OP1
rlabel metal2 4920 960 4932 960 1 LOAD_ACC
rlabel metal2 6024 960 6036 960 1 ACC_INV_Cout
rlabel metal2 6168 960 6180 960 1 INV_REM
rlabel metal2 4200 960 4212 960 1 ACC_Cout
rlabel metal2 1944 960 1956 960 5 INV_OP2
rlabel metal2 2208 960 2220 960 5 DIVH_P
rlabel metal2 2136 960 2148 960 1 LOAD_DIVH
rlabel metal2 7152 960 7164 960 1 RESULT_P
rlabel metal2 8232 960 8244 960 1 RESULT_INV_Cout
rlabel metal2 8376 960 8388 960 1 INV_RESULT
rlabel metal2 6384 960 6396 960 5 LOAD_REM
rlabel metal2 8592 960 8604 960 5 LOAD_QUOT
rlabel metal2 5880 0 5892 0 1 ACC_INV_Cin
rlabel metal2 288 0 300 0 1 nReset
rlabel metal2 264 0 276 0 1 Clock
rlabel metal2 240 0 252 0 1 Test
rlabel metal2 216 0 228 0 1 SDI
rlabel metal2 0 0 200 0 1 Vdd!
rlabel metal2 9360 960 9560 960 5 GND!
rlabel metal2 9360 0 9560 0 1 GND!
rlabel metal2 7128 960 7140 960 5 RESULT_nP_0
rlabel metal1 9570 855 9570 865 7 Quotient
rlabel metal1 9570 902 9570 912 7 Remainder
<< end >>
