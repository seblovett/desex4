magic
tech c035u
timestamp 1387314597
<< metal1 >>
rect 4261 918 5063 928
rect 1861 895 2015 907
rect 4765 896 4919 906
rect 7141 902 9786 912
rect 0 874 4392 884
rect 4406 874 4870 884
rect 4957 874 5111 884
rect 6301 875 6455 885
rect 8509 880 8663 890
rect 0 853 1487 863
rect 1501 852 1967 862
rect 2053 852 2159 862
rect 2245 852 2375 862
rect 3061 854 3191 864
rect 3229 854 3360 864
rect 3781 852 3911 862
rect 3973 852 4055 862
rect 4141 852 5783 862
rect 5797 852 5927 862
rect 5941 852 6407 862
rect 7285 860 7415 870
rect 8005 857 8135 867
rect 8149 857 8615 867
rect 9349 855 9786 865
<< m2contact >>
rect 4247 916 4261 930
rect 5063 916 5077 930
rect 1847 894 1861 908
rect 2015 894 2029 908
rect 4751 894 4765 908
rect 4919 894 4933 908
rect 7127 901 7141 915
rect 4392 872 4406 886
rect 4870 872 4884 886
rect 4943 872 4957 886
rect 5111 872 5125 886
rect 6287 873 6301 887
rect 6455 873 6469 887
rect 8495 878 8509 892
rect 8663 878 8677 892
rect 1487 850 1501 864
rect 1967 850 1981 864
rect 2039 850 2053 864
rect 2159 850 2173 864
rect 2231 850 2245 864
rect 2375 850 2389 864
rect 3047 850 3061 864
rect 3191 850 3205 864
rect 3215 850 3229 864
rect 3360 850 3374 864
rect 3767 850 3781 864
rect 3911 850 3925 864
rect 3959 850 3973 864
rect 4055 850 4069 864
rect 4127 850 4141 864
rect 5783 850 5797 864
rect 5927 850 5941 864
rect 6407 850 6421 864
rect 7271 857 7285 871
rect 7415 858 7429 872
rect 7991 855 8005 869
rect 8135 855 8149 869
rect 8615 855 8629 869
rect 9335 851 9349 865
<< metal2 >>
rect 1536 851 1644 863
rect 1488 847 1500 850
rect 1536 847 1548 851
rect 1632 847 1644 851
rect 1800 847 1812 960
rect 1848 847 1860 894
rect 1944 847 1956 960
rect 1968 847 1980 850
rect 2016 847 2028 894
rect 2040 847 2052 850
rect 2136 847 2148 960
rect 2160 847 2172 850
rect 2208 847 2220 960
rect 2232 847 2244 850
rect 2376 847 2388 850
rect 3000 847 3012 960
rect 3048 847 3060 850
rect 3120 847 3132 960
rect 3144 847 3156 960
rect 3192 847 3204 850
rect 3216 847 3228 850
rect 3360 847 3372 850
rect 3768 847 3780 850
rect 3912 847 3924 850
rect 3960 847 3972 850
rect 4056 847 4068 850
rect 4128 847 4140 850
rect 4248 847 4260 916
rect 4320 847 4332 960
rect 4392 847 4404 872
rect 4440 853 4548 865
rect 4440 847 4452 853
rect 4536 847 4548 853
rect 4704 847 4716 960
rect 4752 847 4764 894
rect 4848 847 4860 960
rect 4872 847 4884 872
rect 4920 847 4932 894
rect 4944 847 4956 872
rect 5040 847 5052 960
rect 5064 847 5076 916
rect 5112 847 5124 872
rect 5136 851 5220 863
rect 5136 847 5148 851
rect 5208 847 5220 851
rect 5256 847 5268 960
rect 5784 847 5796 850
rect 5928 847 5941 850
rect 5976 851 6084 863
rect 5976 847 5988 851
rect 6072 847 6084 851
rect 6240 847 6252 960
rect 6288 847 6300 873
rect 6384 847 6396 960
rect 6408 847 6420 850
rect 6456 847 6468 873
rect 6480 851 6564 863
rect 6480 847 6492 851
rect 6552 847 6564 851
rect 6600 847 6612 960
rect 7128 847 7140 901
rect 7272 847 7284 857
rect 7344 847 7356 960
rect 7368 847 7380 960
rect 7416 847 7428 858
rect 7440 853 7596 865
rect 7440 847 7452 853
rect 7584 847 7596 853
rect 7992 847 8004 855
rect 8136 847 8148 855
rect 8184 854 8292 866
rect 8184 847 8196 854
rect 8280 847 8292 854
rect 8448 847 8460 960
rect 8496 847 8508 878
rect 8592 847 8604 960
rect 8616 847 8628 855
rect 8664 847 8676 878
rect 8688 856 8772 868
rect 8688 847 8700 856
rect 8760 847 8772 856
rect 8808 847 8820 960
rect 9336 847 9348 851
rect 9576 847 9776 960
rect 0 0 200 48
rect 216 0 228 48
rect 240 0 252 48
rect 264 0 276 48
rect 288 0 300 48
rect 1656 0 1668 48
rect 2784 35 2796 48
rect 2928 35 2940 48
rect 2784 23 2940 35
rect 2784 0 2796 23
rect 2952 0 2964 48
rect 3768 0 3780 48
rect 4176 0 4188 48
rect 4560 0 4572 48
rect 5256 0 5268 48
rect 6096 0 6108 48
rect 7992 0 8004 48
rect 8304 0 8316 48
rect 9576 0 9776 48
use leftbuf leftbuf_0
timestamp 1386242881
transform 1 0 0 0 1 48
box 0 0 1464 799
use inv inv_0
timestamp 1386238110
transform 1 0 1464 0 1 48
box 0 0 120 799
use halfadder halfadder_0
timestamp 1386235204
transform 1 0 1584 0 1 48
box 0 0 312 799
use mux2 mux2_0
timestamp 1386235218
transform 1 0 1896 0 1 48
box 0 0 192 799
use mux2 mux2_1
timestamp 1386235218
transform 1 0 2088 0 1 48
box 0 0 192 799
use scandtype scandtype_0
timestamp 1386241841
transform 1 0 2280 0 1 48
box 0 0 624 799
use nor2 nor2_0
timestamp 1386235306
transform 1 0 2904 0 1 48
box 0 0 120 799
use tielow tielow_0
timestamp 1386086605
transform 1 0 3024 0 1 48
box 0 0 48 799
use mux2 mux2_2
timestamp 1386235218
transform 1 0 3072 0 1 48
box 0 0 192 799
use scandtype scandtype_1
timestamp 1386241841
transform 1 0 3264 0 1 48
box 0 0 624 799
use inv inv_4
timestamp 1386238110
transform 1 0 3888 0 1 48
box 0 0 120 799
use fulladder fulladder_0
timestamp 1386234928
transform 1 0 4008 0 1 48
box 0 0 360 799
use inv inv_1
timestamp 1386238110
transform 1 0 4368 0 1 48
box 0 0 120 799
use halfadder halfadder_1
timestamp 1386235204
transform 1 0 4488 0 1 48
box 0 0 312 799
use mux2 mux2_3
timestamp 1386235218
transform 1 0 4800 0 1 48
box 0 0 192 799
use mux2 mux2_4
timestamp 1386235218
transform 1 0 4992 0 1 48
box 0 0 192 799
use scanreg scanreg_2
timestamp 1386241447
transform 1 0 5184 0 1 48
box 0 0 720 799
use inv inv_2
timestamp 1386238110
transform 1 0 5904 0 1 48
box 0 0 120 799
use halfadder halfadder_2
timestamp 1386235204
transform 1 0 6024 0 1 48
box 0 0 312 799
use mux2 mux2_5
timestamp 1386235218
transform 1 0 6336 0 1 48
box 0 0 192 799
use scanreg scanreg_0
timestamp 1386241447
transform 1 0 6528 0 1 48
box 0 0 720 799
use tielow tielow_1
timestamp 1386086605
transform 1 0 7248 0 1 48
box 0 0 48 799
use mux2 mux2_6
timestamp 1386235218
transform 1 0 7296 0 1 48
box 0 0 192 799
use scandtype scandtype_4
timestamp 1386241841
transform 1 0 7488 0 1 48
box 0 0 624 799
use inv inv_3
timestamp 1386238110
transform 1 0 8112 0 1 48
box 0 0 120 799
use halfadder halfadder_3
timestamp 1386235204
transform 1 0 8232 0 1 48
box 0 0 312 799
use mux2 mux2_7
timestamp 1386235218
transform 1 0 8544 0 1 48
box 0 0 192 799
use scanreg scanreg_1
timestamp 1386241447
transform 1 0 8736 0 1 48
box 0 0 720 799
use rightend rightend_0
timestamp 1386235834
transform 1 0 9456 0 1 48
box 0 0 320 799
<< labels >>
rlabel metal1 0 853 0 863 3 Operand2
rlabel metal1 0 874 0 884 4 Operand1
rlabel metal2 1656 0 1668 0 1 OP2_INV_Cin
rlabel metal2 2784 0 2796 0 1 DIVH_1
rlabel metal2 1800 960 1812 960 5 OP2_INV_Cout
rlabel metal2 1944 960 1956 960 5 INV_OP2
rlabel metal2 2208 960 2220 960 5 DIVH_P
rlabel metal2 2136 960 2148 960 1 LOAD_DIVH
rlabel metal2 288 0 300 0 1 nReset
rlabel metal2 264 0 276 0 1 Clock
rlabel metal2 240 0 252 0 1 Test
rlabel metal2 216 0 228 0 1 SDI
rlabel metal2 0 0 200 0 1 Vdd!
rlabel metal2 4560 0 4572 0 1 OP1_INV_Cin
rlabel metal2 3768 0 3780 0 1 DIVL_1
rlabel metal2 4176 0 4188 0 1 ACC_Cin
rlabel metal2 3144 960 3156 960 5 DIVL_P
rlabel metal2 3120 960 3132 960 5 LOAD_DIVL
rlabel metal2 4704 960 4716 960 1 OP1_INV_Cout
rlabel metal2 4848 960 4860 960 5 INV_OP1
rlabel metal2 5040 960 5052 960 1 LOAD_ACC
rlabel metal2 4320 960 4332 960 1 ACC_Cout
rlabel metal2 6240 960 6252 960 1 ACC_INV_Cout
rlabel metal2 6384 960 6396 960 1 INV_REM
rlabel metal2 7368 960 7380 960 1 RESULT_P
rlabel metal2 8448 960 8460 960 1 RESULT_INV_Cout
rlabel metal2 8592 960 8604 960 1 INV_RESULT
rlabel metal2 6600 960 6612 960 5 LOAD_REM
rlabel metal2 8808 960 8820 960 5 LOAD_QUOT
rlabel metal2 7344 960 7356 960 5 RESULT_nP_0
rlabel metal1 9786 855 9786 865 7 Quotient
rlabel metal1 9786 902 9786 912 7 Remainder
rlabel metal2 5256 960 5268 960 5 ACC_LOAD
rlabel metal2 5256 0 5268 0 1 ACC_LOAD
rlabel metal2 2952 0 2964 0 1 DIVH_0_P
rlabel metal2 3000 960 3012 960 5 DIVH_0
rlabel metal2 6096 0 6108 0 1 ACC_INV_Cin
rlabel metal2 8304 0 8316 0 1 RESULT_INV_Cin
rlabel metal2 7992 0 8004 0 1 RESULT_1
rlabel metal2 9576 0 9776 0 1 GND!
rlabel metal2 9576 960 9776 960 5 GND!
<< end >>
